package parameters_pkg;
parameter int DATA_WIDTH = 448;
// p = 2^448 - 2^224 - 1
parameter logic [DATA_WIDTH-1:0] MODULUS = 448'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
parameter logic [DATA_WIDTH-1:0] MODULUS_INV = 448'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000001;
// R = 2^448
parameter logic [DATA_WIDTH:0] R = 449'h10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
parameter logic [DATA_WIDTH-1:0] R_MOD_P = 448'h100000000000000000000000000000000000000000000000000000001;
parameter logic [DATA_WIDTH-1:0] R_INV = 448'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000001;
parameter logic [DATA_WIDTH-1:0] R2_MOD_P = 448'h0000000000000000000000000000000000000000000000000000000300000000000000000000000000000000000000000000000000000002;

// d = -39081
// D = d*R Montgomery representation
parameter logic [DATA_WIDTH-1:0] D = 448'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6755FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6756;
endpackage